module main

import vjvm

fn main() {
}
